`ifndef TLB_PARAMS_SVH
`define TLB_PARAMS_SVH



`endif