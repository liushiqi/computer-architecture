

module pipeline;