package axi_params;
typedef logic [31:0] AXIData;
endpackage;

module cpu_axi_interface (
  input clock,
  input reset_,
  input instruction_ram_request,
  input instruction_ram_write,
  input [1:0] instruction_ram_size,
  input axi_params::AXIData instruction_ram_address,
  input axi_params::AXIData instruction_ram_write_data,
  output axi_params::AXIData instruction_ram_read_data,
  output instruction_ram_address_ready,
  output instruction_ram_data_ready,
  input data_ram_request,
  input data_ram_write,
  input [1:0] data_ram_size,
  input axi_params::AXIData data_ram_address,
  input axi_params::AXIData data_ram_write_data,
  output axi_params::AXIData data_ram_read_data,
  output data_ram_address_ready,
  output data_ram_data_ready,
  output [3:0] axi_read_address_id,
  output axi_params::AXIData axi_read_address,
  output [7:0] axi_read_address_length,
  output [2:0] axi_read_address_size,
  output [1:0] axi_read_address_burst,
  output [1:0] axi_read_address_lock,
  output [3:0] axi_read_address_cache,
  output [2:0] axi_read_address_protection,
  output axi_read_address_valid,
  input axi_read_address_ready,
  input [3:0] axi_read_data_id,
  input axi_params::AXIData axi_read_data,
  input [1:0] axi_read_data_response,
  input axi_read_data_last,
  input axi_read_data_valid,
  output axi_read_data_ready,
  output [3:0] axi_write_address_id,
  output axi_params::AXIData axi_write_address,
  output [7:0] axi_write_address_length,
  output [2:0] axi_write_address_size,
  output [1:0] axi_write_address_burst,
  output [1:0] axi_write_address_lock,
  output [3:0] axi_write_address_cache,
  output [2:0] axi_write_address_protection,
  output axi_write_address_valid,
  input axi_write_address_ready,
  output [3:0] axi_write_data_id,
  output axi_params::AXIData axi_write_data,
  output [3:0] axi_write_data_strobe,
  output axi_write_data_last,
  output axi_write_data_valid,
  input axi_write_data_ready,
  input [3:0] axi_write_responce_id,
  input [1:0] axi_write_responce,
  input axi_write_responce_valid,
  output axi_write_responce_ready
);
  import axi_params::*;
  wire reset;
  assign reset = ~reset_;
endmodule